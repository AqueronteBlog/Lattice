/* Verilog model created from schematic LED_Blinky.sch -- Dec 25, 2018 23:15 */

module LED_Blinky;




endmodule // LED_Blinky
